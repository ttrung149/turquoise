signal logic : std_logic;
signal logic_vector_1, logic_vector_2 : std_logic_vector(3 downto 0);
signal int_1, int_2, int_3 : integer := 42;
signal u : unsigned(3 downto 0);
signal s : signed(3 downto 0);
signal a, b, c : string := "hello world";